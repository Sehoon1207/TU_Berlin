entity BLACK_BOX is
    port(A,B : in std_logic;
         C   : out std_logic);
end entity BLACK_BOX;